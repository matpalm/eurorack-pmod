po2_network.sv