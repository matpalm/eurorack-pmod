qb_network.sv